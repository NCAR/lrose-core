netcdf KRAX {
dimensions:
	Time = UNLIMITED ;
	numSystems = 1 ;
	long_string = 80 ;
variables:
	int volume_start_time ;
		volume_start_time:long_name = "Unix Date/Time value for volume start time" ;
		volume_start_time:units = "seconds since 1970-01-01 00:00 UTC" ;
	int base_time ;
		base_time:long_name = "Unix Date/Time value for first record" ;
		base_time:units = "seconds since 1970-01-01 00:00 UTC" ;
		base_time:missing_value = 0 ;
		base_time:_FillValue = 0 ;
	float Fixed_Angle ;
		Fixed_Angle:long_name = "Targeted fixed angle for this scan" ;
		Fixed_Angle:units = "degrees" ;
		Fixed_Angle:missing_value = -32768.f ;
		Fixed_Angle:_FillValue = -32768.f ;
	float Nyquist_Velocity ;
		Nyquist_Velocity:long_name = "Effective unambigous velocity" ;
		Nyquist_Velocity:units = "meters/second" ;
		Nyquist_Velocity:missing_value = -32768.f ;
		Nyquist_Velocity:_FillValue = -32768.f ;
	float Unambiguous_Range ;
		Unambiguous_Range:long_name = "Effective unambigous range" ;
		Unambiguous_Range:units = "kilometers" ;
		Unambiguous_Range:missing_value = -32768.f ;
		Unambiguous_Range:_FillValue = -32768.f ;
	double Latitude ;
		Latitude:long_name = "Latitude of the instrument" ;
		Latitude:units = "degrees_north" ;
		Latitude:valid_range = -90.f, 90.f ;
		Latitude:missing_value = -32768. ;
		Latitude:_FillValue = -32768. ;
	double Longitude ;
		Longitude:long_name = "Longitude of the instrument" ;
		Longitude:units = "degrees_east" ;
		Longitude:valid_range = -360.f, 360.f ;
		Longitude:missing_value = -32768. ;
		Longitude:_FillValue = -32768. ;
	double Altitude ;
		Altitude:long_name = "Altitude in meters (asl) of the instrument" ;
		Altitude:units = "meters" ;
		Altitude:valid_range = -10000., 90000. ;
		Altitude:missing_value = -32768. ;
		Altitude:_FillValue = -32768. ;
	float Radar_Constant(numSystems) ;
		Radar_Constant:long_name = "Radar constant" ;
		Radar_Constant:units = "???" ;
		Radar_Constant:missing_value = -32768.f ;
		Radar_Constant:_FillValue = -32768.f ;
	float rcvr_gain(numSystems) ;
		rcvr_gain:long_name = "Receiver Gain" ;
		rcvr_gain:Comment = "Most entries are 2 dimension arrays one for each polarity" ;
		rcvr_gain:units = "db" ;
		rcvr_gain:missing_value = -32768.f ;
		rcvr_gain:_FillValue = -32768.f ;
	float ant_gain(numSystems) ;
		ant_gain:long_name = "Antenna Gain" ;
		ant_gain:units = "db" ;
		ant_gain:missing_value = -32768.f ;
		ant_gain:_FillValue = -32768.f ;
	float sys_gain(numSystems) ;
		sys_gain:long_name = "System Gain" ;
		sys_gain:units = "db" ;
		sys_gain:missing_value = -32768.f ;
		sys_gain:_FillValue = -32768.f ;
	float bm_width(numSystems) ;
		bm_width:long_name = "Beam Width" ;
		bm_width:units = "degrees" ;
		bm_width:missing_value = -32768.f ;
		bm_width:_FillValue = -32768.f ;
	float pulse_width(numSystems) ;
		pulse_width:long_name = "Pulse Width" ;
		pulse_width:units = "seconds" ;
		pulse_width:missing_value = -32768.f ;
		pulse_width:_FillValue = -32768.f ;
	float band_width(numSystems) ;
		band_width:long_name = "Band Width" ;
		band_width:units = "hertz" ;
		band_width:missing_value = -32768.f ;
		band_width:_FillValue = -32768.f ;
	float peak_pwr(numSystems) ;
		peak_pwr:long_name = "Peak Power" ;
		peak_pwr:units = "watts" ;
		peak_pwr:missing_value = -32768.f ;
		peak_pwr:_FillValue = -32768.f ;
	float xmtr_pwr(numSystems) ;
		xmtr_pwr:long_name = "Transmitter Power" ;
		xmtr_pwr:units = "dBm" ;
		xmtr_pwr:missing_value = -32768.f ;
		xmtr_pwr:_FillValue = -32768.f ;
	float noise_pwr(numSystems) ;
		noise_pwr:long_name = "Noise Power" ;
		noise_pwr:units = "dBm" ;
		noise_pwr:missing_value = -32768.f ;
		noise_pwr:_FillValue = -32768.f ;
	float tst_pls_pwr(numSystems) ;
		tst_pls_pwr:long_name = "Test Pulse Power" ;
		tst_pls_pwr:units = "dBm" ;
		tst_pls_pwr:missing_value = -32768.f ;
		tst_pls_pwr:_FillValue = -32768.f ;
	float tst_pls_rng0(numSystems) ;
		tst_pls_rng0:long_name = "Range to start of test pulse" ;
		tst_pls_rng0:units = "meters" ;
		tst_pls_rng0:missing_value = -32768.f ;
		tst_pls_rng0:_FillValue = -32768.f ;
	float tst_pls_rng1(numSystems) ;
		tst_pls_rng1:long_name = "Range to end of test pulse" ;
		tst_pls_rng1:units = "meters" ;
		tst_pls_rng1:missing_value = -32768.f ;
		tst_pls_rng1:_FillValue = -32768.f ;
	float Wavelength(numSystems) ;
		Wavelength:long_name = "System wavelength" ;
		Wavelength:units = "meters" ;
		Wavelength:missing_value = -32768.f ;
		Wavelength:_FillValue = -32768.f ;
	float PRF(numSystems) ;
		PRF:long_name = "System pulse repetition frequence" ;
		PRF:units = "pulses/sec" ;
		PRF:missing_value = -32768.f ;
		PRF:_FillValue = -32768.f ;
	float sur_PRF(numSystems) ;
		sur_PRF:long_name = "PRF for surveillance sweep if combined" ;
		sur_PRF:units = "pulses/sec" ;
		sur_PRF:missing_value = -32768.f ;
		sur_PRF:_FillValue = -32768.f ;
	float dbz0(numSystems) ;
		dbz0:long_name = "Scaling constant used by the signal processor to calculate reflectivity" ;
		dbz0:units = "dB" ;
		dbz0:missing_value = -32768.f ;
		dbz0:_FillValue = -32768.f ;
	float horiz_noise(numSystems) ;
		horiz_noise:long_name = " Noise level horizontal channel" ;
		horiz_noise:units = "dBm" ;
		horiz_noise:missing_value = -32768.f ;
		horiz_noise:_FillValue = -32768.f ;
	float vert_noise(numSystems) ;
		vert_noise:long_name = " Noise level vertical channel" ;
		vert_noise:units = "dBm" ;
		vert_noise:missing_value = -32768.f ;
		vert_noise:_FillValue = -32768.f ;
	float channel_config(numSystems) ;
		channel_config:long_name = "Channel Configuration" ;
		channel_config:units = "coded" ;
		channel_config:missing_value = -32768.f ;
		channel_config:_FillValue = -32768.f ;
	float waveform_type(numSystems) ;
		waveform_type:long_name = "Waveform Type" ;
		waveform_type:units = "coded" ;
		waveform_type:missing_value = -32768.f ;
		waveform_type:_FillValue = -32768.f ;
	float super_res_control(numSystems) ;
		super_res_control:long_name = "Super Resolution Control" ;
		super_res_control:units = "coded" ;
		super_res_control:missing_value = -32768.f ;
		super_res_control:_FillValue = -32768.f ;
	float sur_prf_num(numSystems) ;
		sur_prf_num:long_name = "Surveillance PRF Number" ;
		sur_prf_num:units = "n/a" ;
		sur_prf_num:missing_value = -32768.f ;
		sur_prf_num:_FillValue = -32768.f ;
	float sur_prf_pulse_count(numSystems) ;
		sur_prf_pulse_count:long_name = "Surveillance PRF pulse count per radial" ;
		sur_prf_pulse_count:units = "n/a" ;
		sur_prf_pulse_count:missing_value = -32768.f ;
		sur_prf_pulse_count:_FillValue = -32768.f ;
	float dop_prf_num(numSystems) ;
		dop_prf_num:long_name = "Doppler PRF Number" ;
		dop_prf_num:units = "n/a" ;
		dop_prf_num:missing_value = -32768.f ;
		dop_prf_num:_FillValue = -32768.f ;
	float dop_prf_pulse_count(numSystems) ;
		dop_prf_pulse_count:long_name = "Doppler PRF pulse count per radial" ;
		dop_prf_pulse_count:units = "n/a" ;
		dop_prf_pulse_count:missing_value = -32768.f ;
		dop_prf_pulse_count:_FillValue = -32768.f ;
	float azimuth_rate(numSystems) ;
		azimuth_rate:long_name = "Azimuth scan rate" ;
		azimuth_rate:units = "deg/s" ;
		azimuth_rate:missing_value = -32768.f ;
		azimuth_rate:_FillValue = -32768.f ;
	int RDA_build_num(numSystems) ;
		RDA_build_num:long_name = "RDA major and minor build number" ;
		RDA_build_num:units = "n/a" ;
		RDA_build_num:missing_value = 0 ;
		RDA_build_num:_FillValue = 0 ;
	double time_offset(Time) ;
		time_offset:long_name = "time offset of the current record from base_time" ;
		time_offset:units = "seconds" ;
		time_offset:missing = -32768. ;
		time_offset:_FillValue = -32768. ;
	float Azimuth(Time) ;
		Azimuth:long_name = "Earth relative azimuth of the ray" ;
		Azimuth:Comment = "Degrees clockwise from true North" ;
		Azimuth:units = "degrees" ;
		Azimuth:valid_range = -360.f, 360.f ;
		Azimuth:missing_value = -32768.f ;
		Azimuth:_FillValue = -32768.f ;
	float Elevation(Time) ;
		Elevation:long_name = "Earth relative elevation of the ray" ;
		Elevation:Comment = "Degrees from earth tangent towards zenith" ;
		Elevation:units = "degrees" ;
		Elevation:valid_range = -360.f, 360.f ;
		Elevation:missing_value = -32768.f ;
		Elevation:_FillValue = -32768.f ;
	float clip_range(Time) ;
		clip_range:long_name = "Range of last usefull cell" ;
		clip_range:units = "meters" ;
		clip_range:missing_value = -32768.f ;
		clip_range:_FillValue = -32768.f ;

}
